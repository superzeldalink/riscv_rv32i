// `ifdef SIMULATION
parameter IMEM_DEPTH = 8192;
parameter DMEM_DEPTH = 2048;
// `else
// parameter IMEM_DEPTH = 1024;
// parameter DMEM_DEPTH = 128;
// `endif
